LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
use ieee.numeric_std.all;

entity my_base_tempo is
	Generic ( DATA_SIZE : natural := 8;
				 BT_RAPIDO : natural := 25000000);
    port(
        clk      :   in std_logic;
        sw_in : in std_logic;
        enable : in std_logic;
		  
		  reset : in std_logic;
		  readEnable : in std_logic;
		  writeEnable : in std_logic;
		  
		  ledRapido : out std_logic;
		 
        saida_clk :   out std_logic_vector(DATA_SIZE-1 downto 0)
        );
end entity;

architecture divInteiro of my_base_tempo is
    signal tick : std_logic := '0';
    signal divisor : natural := 50000000;
    signal contador : integer range 0 to 100000000 := 0;
begin
    -- sw seleciona o divisor
	 divisor <= 50000000 when sw_in='0' else BT_RAPIDO;
	 ledRapido <= sw_in;
   process(clk)
    begin
        if rising_edge(clk) then
				if (reset='1') then
					contador <= 0;
            -- contador e comparador
            elsif contador >= divisor then
--                contador <= 0;
                tick <= '1';
            else
                contador <= contador + 1;
					 tick <= '0';
            end if;
        end if;
	end process;
   -- saida do clock em 8 bits quando enable, no contrário saida é impedância
	saida_clk <= ("0000000" & tick) when (enable='1' AND readEnable='1') else "ZZZZZZZZ";
end architecture divInteiro;