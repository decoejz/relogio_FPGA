
library IEEE;
use ieee.std_logic_1164.all;

entity my_base_tempo is
    port
    (
       A : in std_logic
    );
end entity;

architecture base_tempoArc of my_base_tempo is


begin

	
end architecture;