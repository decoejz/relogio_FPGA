
library IEEE;
use ieee.std_logic_1164.all;

entity relogio is
    port
    (
       A : in std_logic
    );
end entity;

architecture relogioArc of relogio is


begin
    
end architecture;