
library IEEE;
use ieee.std_logic_1164.all;

entity my_processador is
    port
    (
       A : in std_logic
    );
end entity;

architecture processadorArc of my_processador is


begin
    
end architecture;