
library IEEE;
use ieee.std_logic_1164.all;

entity my_pc is
    port
    (
       A : in std_logic
    );
end entity;

architecture pcArc of my_pc is


begin

	
end architecture;