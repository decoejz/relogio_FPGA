
library IEEE;
use ieee.std_logic_1164.all;

entity my_flip_flop is
    port
    (
       A : in std_logic
    );
end entity;

architecture flip_flopArc of my_flip_flop is


begin

	
end architecture;