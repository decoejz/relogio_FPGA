
library IEEE;
use ieee.std_logic_1164.all;

entity my_tristate is
    port
    (
       A : in std_logic
    );
end entity;

architecture tristateArc of my_tristate is


begin

	
end architecture;